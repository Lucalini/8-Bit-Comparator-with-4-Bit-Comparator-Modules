`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/01/2023 05:17:13 PM
// Design Name: 
// Module Name: Fourbitcomparator
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Fourbitcomparator(
    input [3:0] a,
    input [3:0] b,
    output eq,
    output lt,
    output gt
    );
endmodule
